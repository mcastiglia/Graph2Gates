module main(a,b,s,cout);
input [31:0] a,b;
output [31:0] s;
output cout;
wire g0_0,g22_22,p26_26,c11,c8,p23_23,c24,c27,p10_10,g13_0,p28_28,p20_20,p30_30,c0,c26,p4_4,g11_11,c29,g23_0,g22_0,p19_19,g16_16,g1_1,c13,p31_31,g27_0,p15_15,g15_0,g28_0,p29_29,c19,g14_0,c3,g6_6,p5_5,g21_0,g21_21,g25_0,g20_0,c30,p16_16,p2_2,g8_0,c2,g16_0,c6,c10,c25,g17_0,p17_17,g24_24,g4_0,c20,g24_0,g12_0,g28_28,g10_0,p22_22,g5_5,c7,c12,p25_25,g9_0,g2_0,c31,g29_0,p18_18,g26_26,c15,g25_25,p7_7,g6_0,g3_3,g17_17,p14_14,p9_9,c18,p21_21,g18_18,g26_0,g14_14,g8_8,p6_6,c9,p0_0,c22,c16,p27_27,p13_13,g2_2,p12_12,c28,c5,g7_0,g29_29,g9_9,c1,g10_10,c14,p8_8,p1_1,g23_23,g1_0,c4,g13_13,g27_27,c21,g15_15,g18_0,g7_7,g19_19,p11_11,p3_3,c17,g5_0,g12_12,g19_0,g30_0,g30_30,g31_31,c23,g20_20,p24_24,g11_0,g4_4,g3_0;

assign p0_0 = a[0] ^ b[0];
assign g0_0 = a[0] & b[0];
assign p1_1 = a[1] ^ b[1];
assign g1_1 = a[1] & b[1];
assign p2_2 = a[2] ^ b[2];
assign g2_2 = a[2] & b[2];
assign p3_3 = a[3] ^ b[3];
assign g3_3 = a[3] & b[3];
assign p4_4 = a[4] ^ b[4];
assign g4_4 = a[4] & b[4];
assign p5_5 = a[5] ^ b[5];
assign g5_5 = a[5] & b[5];
assign p6_6 = a[6] ^ b[6];
assign g6_6 = a[6] & b[6];
assign p7_7 = a[7] ^ b[7];
assign g7_7 = a[7] & b[7];
assign p8_8 = a[8] ^ b[8];
assign g8_8 = a[8] & b[8];
assign p9_9 = a[9] ^ b[9];
assign g9_9 = a[9] & b[9];
assign p10_10 = a[10] ^ b[10];
assign g10_10 = a[10] & b[10];
assign p11_11 = a[11] ^ b[11];
assign g11_11 = a[11] & b[11];
assign p12_12 = a[12] ^ b[12];
assign g12_12 = a[12] & b[12];
assign p13_13 = a[13] ^ b[13];
assign g13_13 = a[13] & b[13];
assign p14_14 = a[14] ^ b[14];
assign g14_14 = a[14] & b[14];
assign p15_15 = a[15] ^ b[15];
assign g15_15 = a[15] & b[15];
assign p16_16 = a[16] ^ b[16];
assign g16_16 = a[16] & b[16];
assign p17_17 = a[17] ^ b[17];
assign g17_17 = a[17] & b[17];
assign p18_18 = a[18] ^ b[18];
assign g18_18 = a[18] & b[18];
assign p19_19 = a[19] ^ b[19];
assign g19_19 = a[19] & b[19];
assign p20_20 = a[20] ^ b[20];
assign g20_20 = a[20] & b[20];
assign p21_21 = a[21] ^ b[21];
assign g21_21 = a[21] & b[21];
assign p22_22 = a[22] ^ b[22];
assign g22_22 = a[22] & b[22];
assign p23_23 = a[23] ^ b[23];
assign g23_23 = a[23] & b[23];
assign p24_24 = a[24] ^ b[24];
assign g24_24 = a[24] & b[24];
assign p25_25 = a[25] ^ b[25];
assign g25_25 = a[25] & b[25];
assign p26_26 = a[26] ^ b[26];
assign g26_26 = a[26] & b[26];
assign p27_27 = a[27] ^ b[27];
assign g27_27 = a[27] & b[27];
assign p28_28 = a[28] ^ b[28];
assign g28_28 = a[28] & b[28];
assign p29_29 = a[29] ^ b[29];
assign g29_29 = a[29] & b[29];
assign p30_30 = a[30] ^ b[30];
assign g30_30 = a[30] & b[30];
assign p31_31 = a[31] ^ b[31];
assign g31_31 = a[31] & b[31];
assign g1_0 = c1;
assign g2_0 = c2;
assign g3_0 = c3;
assign g4_0 = c4;
assign g5_0 = c5;
assign g6_0 = c6;
assign g7_0 = c7;
assign g8_0 = c8;
assign g9_0 = c9;
assign g10_0 = c10;
assign g11_0 = c11;
assign g12_0 = c12;
assign g13_0 = c13;
assign g14_0 = c14;
assign g15_0 = c15;
assign g16_0 = c16;
assign g17_0 = c17;
assign g18_0 = c18;
assign g19_0 = c19;
assign g20_0 = c20;
assign g21_0 = c21;
assign g22_0 = c22;
assign g23_0 = c23;
assign g24_0 = c24;
assign g25_0 = c25;
assign g26_0 = c26;
assign g27_0 = c27;
assign g28_0 = c28;
assign g29_0 = c29;
assign g30_0 = c30;
assign g31_0 = c31;
GREY grey31(g31_31, p31_31, g30_0, c31);
GREY grey30(g30_30, p30_30, g29_0, c30);
GREY grey29(g29_29, p29_29, g28_0, c29);
GREY grey28(g28_28, p28_28, g27_0, c28);
GREY grey27(g27_27, p27_27, g26_0, c27);
GREY grey26(g26_26, p26_26, g25_0, c26);
GREY grey25(g25_25, p25_25, g24_0, c25);
GREY grey24(g24_24, p24_24, g23_0, c24);
GREY grey23(g23_23, p23_23, g22_0, c23);
GREY grey22(g22_22, p22_22, g21_0, c22);
GREY grey21(g21_21, p21_21, g20_0, c21);
GREY grey20(g20_20, p20_20, g19_0, c20);
GREY grey19(g19_19, p19_19, g18_0, c19);
GREY grey18(g18_18, p18_18, g17_0, c18);
GREY grey17(g17_17, p17_17, g16_0, c17);
GREY grey16(g16_16, p16_16, g15_0, c16);
GREY grey15(g15_15, p15_15, g14_0, c15);
GREY grey14(g14_14, p14_14, g13_0, c14);
GREY grey13(g13_13, p13_13, g12_0, c13);
GREY grey12(g12_12, p12_12, g11_0, c12);
GREY grey11(g11_11, p11_11, g10_0, c11);
GREY grey10(g10_10, p10_10, g9_0, c10);
GREY grey9(g9_9, p9_9, g8_0, c9);
GREY grey8(g8_8, p8_8, g7_0, c8);
GREY grey7(g7_7, p7_7, g6_0, c7);
GREY grey6(g6_6, p6_6, g5_0, c6);
GREY grey5(g5_5, p5_5, g4_0, c5);
GREY grey4(g4_4, p4_4, g3_0, c4);
GREY grey3(g3_3, p3_3, g2_0, c3);
GREY grey2(g2_2, p2_2, g1_0, c2);
GREY grey1(g1_1, p1_1, g0_0, c1);
assign s[0] = a[0] ^ b[0];
assign c0 = g0_0;
assign cout = c31;
assign s[1] = p1_1 ^ c0;
assign s[2] = p2_2 ^ c1;
assign s[3] = p3_3 ^ c2;
assign s[4] = p4_4 ^ c3;
assign s[5] = p5_5 ^ c4;
assign s[6] = p6_6 ^ c5;
assign s[7] = p7_7 ^ c6;
assign s[8] = p8_8 ^ c7;
assign s[9] = p9_9 ^ c8;
assign s[10] = p10_10 ^ c9;
assign s[11] = p11_11 ^ c10;
assign s[12] = p12_12 ^ c11;
assign s[13] = p13_13 ^ c12;
assign s[14] = p14_14 ^ c13;
assign s[15] = p15_15 ^ c14;
assign s[16] = p16_16 ^ c15;
assign s[17] = p17_17 ^ c16;
assign s[18] = p18_18 ^ c17;
assign s[19] = p19_19 ^ c18;
assign s[20] = p20_20 ^ c19;
assign s[21] = p21_21 ^ c20;
assign s[22] = p22_22 ^ c21;
assign s[23] = p23_23 ^ c22;
assign s[24] = p24_24 ^ c23;
assign s[25] = p25_25 ^ c24;
assign s[26] = p26_26 ^ c25;
assign s[27] = p27_27 ^ c26;
assign s[28] = p28_28 ^ c27;
assign s[29] = p29_29 ^ c28;
assign s[30] = p30_30 ^ c29;
assign s[31] = p31_31 ^ c30;
endmodule

module GREY(gik, pik, gkj, gij);
input gik, pik, gkj;
output gij;
assign gij = gik | (pik & gkj);
endmodule

module BLACK(gik, pik, gkj, pkj, gij, pij);
input gik, pik, gkj, pkj;
output gij, pij;
assign pij = pik & pkj;
assign gij = gik | (pik & gkj);
endmodule

